package sfifo_sequence_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;
	
	// importing packages : agent,
	import sfifo_agent_pkg::*;
	
	// include Sequence file:
	`include "sfifo_sequence.svh"
	
endpackage