package sfifo_test_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	
	// import sfifo_pkg::*;
	import sfifo_sequence_pkg::*;
	import sfifo_agent_pkg::*;
	import sfifo_environment_pkg::*;
	
	`include "sfifo_test.svh"
endpackage